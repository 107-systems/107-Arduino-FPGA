---------------------------------------------------------------
-- Viper Quadcopter MKR VIDOR 4000 FPGA Code
-- (C) Alexander Entinger, MSc / LXRobotics GmbH
-- GNU LGPL V3.0
---------------------------------------------------------------

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package RgbLedDefs is

  type aRgbLedColour is (Black, White, Red, Green, Blue, Yellow, Cyan, Magenta);

end RgbLedDefs;
